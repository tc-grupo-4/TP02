*#D:\DATA\MY CIRCUITS\LM833\LM833.CIR SETUP1
*#SAVE V(1) V(4) @VCC[I] @VCC[P] V(2) @R1[I] @R1[P] @R2[I]
*#SAVE @R2[P] V(5) @VEE[I] @VEE[P] @RLOAD[I] @RLOAD[P] V(3)
*#ALIAS VOUT  V(2)
*#VIEW  TRAN VOUT -10V 10V
*#ALIAS VIN  V(3)
*#VIEW  TRAN VIN -10V 10V
*#.TRAN 5N 50U
*#.PRINT  TRAN VOUT
*#.PRINT  TRAN VIN
X1 0 1 4 5 2 LM833#0
*{  }
.SUBCKT LM833#0 1 2 3 4 5
*
C1   11 12 3.501E-12
C2    6  7 10.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 27.96E6
+ -30E6 30E6 30E6 -30E6
GA    6  0 11 12 565.5E-6
GCM   0  6 10 99 5.655E-9
ISS  10  4 DC 70.00E-6
HLIM 90  0 VLIM 1K
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1   3 11 1.768E3
RD2   3 12 1.768E3
RO1   8  5 10
RO2   7 99 20
RP    3  4 29.03E3
RSS  10 99 2.857E6
VB    9  0 DC 0
VC    3 53 DC .9
VE   54  4 DC .4
VLIM  7  8 DC 0
VLP  91  0 DC 30
VLN   0 92 DC 30
.MODEL DX D(IS=800.0E-18)
.MODEL JX NJF(IS=150.0E-9 BETA=4.568E-3
+ VTO=-1)
.ENDS
X2 3 0 SINE#0
*{ AMPLITUDE=3.0V FREQ=100000 }
.SUBCKT SINE#0 1 2
*PARAMETERS:
* OFFSET DC VOLTAGE OFFSET IN VOLTS
* AMP AMPLITUDE IN VOLTS
* FREQ FREQUENCY IN HZ
* DELAY TIME DELAY IN SECONDS
* DAMP DAMPING FACTOR (SEE SIN SOURCE FOR DEFINITION)
V1 1 2 SIN 0 3.0000  100.000K 0 0
R1 1 2 1MEG
.ENDS
VCC 4 0 DC=15.0V
R1 3 1 1.5K
R2 1 2 4.5K
VEE 5 0 DC=-15.0V
RLOAD 2 0 500
.END
